`ifndef SIGNAL_CONNECT__SV
`define SIGNAL_CONNECT__SV

logic		    clk;   
logic 		    rst;   
wire 		    sda;
logic		    scl;   
logic [7:0]	    myReg0;   

logic		    rst_n;
initial 
begin

end


`endif
