`ifndef AD_CHN_IIC_INTERFACE__SV
`define AD_CHN_IIC_INTERFACE__SV

interface ad_chn_iic_interface (input clk, input rst_n);

    logic iic_scl;
    logic iic_sda;

endinterface

`endif
 
